module main;
	initial
	begin
		$display("V is for Verilog");
		$finish;
	end
endmodule

